-- in: from_dout (8 bits)
-- out: to_m_in (18 bits)
